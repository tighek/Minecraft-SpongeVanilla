docker build -t tighek/Minecraft-SpongeVanilla:420B343 .
docker rmi tighek/Minecraft-SpongeVanilla:latest
docker tag tighek/Minecraft-SpongeVanilla:420B343 tighek/Minecraft-SpongeVanilla:latest

